//im dk`
