// im KONDAACHARYULU DITTAKAVI this is a dummy file 
// im creating for practice purpose 
// im a verification engineer
