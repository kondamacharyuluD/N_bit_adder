// im KONDAACHARYULU DITTAKAVI this is a dummy file
