// im KONDAACHARYULU DITTAKAVI this is a dummy fil
// e
