//this is the third practice file
//
//
//
